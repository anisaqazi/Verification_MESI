import master_uvc_pkg::*;
`include "uvm_macros.svh"
import uvm_pkg::*;

`include "mesi_isc_subscriber.sv"
`include "mesi_tb_env.sv"
`include "tests/test_list.sv"
